library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tb_cpu is
generic (
    N : integer := 8                                     -- Number of bit
);
end tb_cpu;

architecture rtl of tb_cpu is
begin

end rtl;
